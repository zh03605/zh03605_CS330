library verilog;
use verilog.vl_types.all;
entity tb2 is
end tb2;
