library verilog;
use verilog.vl_types.all;
entity TB2 is
end TB2;
