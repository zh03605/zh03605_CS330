library verilog;
use verilog.vl_types.all;
entity tb3 is
end tb3;
