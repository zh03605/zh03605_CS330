library verilog;
use verilog.vl_types.all;
entity TB1 is
end TB1;
